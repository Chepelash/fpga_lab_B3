module sorting_tb;



endmodule
